
class eth_pkt_mon;

